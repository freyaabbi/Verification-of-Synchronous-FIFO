`include "generator.sv"
`include "driver.sv"
`include "monitor.sv"
`include "scoreboard.sv"
class environment;
  mailbox gen2drv;
  mailbox mon2scb;
  mailbox gen2scb;

  generator gen;
  driver drv;
  monitor mon;
  scoreboard scb;

  virtual fifo_intf vif;
  event done;
  event clk;

  function new(virtual fifo_intf vif);
    this.vif = vif;
    gen2drv = new();
    mon2scb = new();
    gen2scb = new();
    gen = new(gen2drv, gen2scb);
    drv = new(gen2drv, vif);
    mon = new(mon2scb, vif);
    scb = new(mon2scb, gen2scb);
    gen.done = done;
    scb.done = done;
  endfunction

  task run();
    fork
      gen.main();
      drv.main();
      mon.main();
      scb.main();
    join
  endtask
endclass
